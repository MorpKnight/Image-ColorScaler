LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY DECODER IS
    PORT (
        PROGRAM_COUNTER : IN INTEGER;
        INSTRUCTION : IN STD_LOGIC_VECTOR(49 DOWNTO 0);
        OPCODE : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
    );
END ENTITY DECODER;

ARCHITECTURE DECODE OF DECODER IS

BEGIN

    DEC : PROCESS (PROGRAM_COUNTER, INSTRUCTION)
    BEGIN
        OPCODE <= INSTRUCTION(49 DOWNTO 44);
    END PROCESS DEC;

END ARCHITECTURE DECODE;