LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY DECODER IS
    PORT (
        PROGRAM_COUNTER : IN INTEGER;
        INSTRUCTION : IN STD_LOGIC_VECTOR(0 TO 49);
        OPCODE : OUT STD_LOGIC_VECTOR(0 TO 5)
    );
END ENTITY DECODER;

ARCHITECTURE DECODE OF DECODER IS

BEGIN

    DEC : PROCESS (PROGRAM_COUNTER, INSTRUCTION)
    BEGIN
        OPCODE <= INSTRUCTION(0 TO 5);
    END PROCESS DEC;

END ARCHITECTURE DECODE;