library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SCALER is
    port (
        WIDTH, HEIGHT : in integer;
    );
end entity SCALER;

architecture IMAGESCALLER of SCALER is
    
begin
    
    
    
end architecture IMAGESCALLER;